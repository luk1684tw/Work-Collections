//Subject:     Architecture project 2 - Adder
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//Writer:      
//----------------------------------------------
//Date:        
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------

module Adder(
    src1_i,
	src2_i,
	sum_o
	);
     
	//I/O ports
	input  signed [32-1:0]  src1_i;
	input  signed [32-1:0]	src2_i;
	output signed [32-1:0]	 sum_o;

	//Internal Signals
	wire    [32-1:0]	 sum_o;
//Parameter
    
//Main function
	assign sum_o = src1_i + src2_i;
endmodule